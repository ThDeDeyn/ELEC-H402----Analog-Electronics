** Profile: "SCHEMATIC1-TRAN"  [ D:\PM\Documents PM\Cours\_Analogique\ELEC-H-402 2013-2014\Labos\Labo4 MOS2\Ampli Drain Commun\amplidraincommun-pspicefiles\schematic1\tran.sim ] 

** Creating circuit file "TRAN.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "D:/pm/Documents PM/Cours/_Analogique/ELEC-H-402 2011-2012/Labos/Labo H402 PSpice Lib/small_signal.lib" 
* From [PSPICE NETLIST] section of C:\Program Files\CAO\OrCAD_16.3_Demo\tools\PSpice\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 10m 0 10u 
.FOUR 1k 10 V([Vout]) 
.STEP LIN PARAM DeltaVin 1 2.5 .5 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
