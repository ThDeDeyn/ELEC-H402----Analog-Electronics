** Profile: "SCHEMATIC1-AC"  [ D:\PM\Documents PM\Cours\_Analogique\ELEC-H-402 2013-2014\Labos\Labo4 MOS2\Ampli Drain Commun\amplidraincommun-pspicefiles\schematic1\ac.sim ] 

** Creating circuit file "AC.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "D:/pm/Documents PM/Cours/_Analogique/ELEC-H-402 2011-2012/Labos/Labo H402 PSpice Lib/small_signal.lib" 
* From [PSPICE NETLIST] section of C:\Program Files\CAO\OrCAD_16.3_Demo\tools\PSpice\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 5 1Hz 1GHz
.STEP PARAM RLval LIST 100Meg,20 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
