** Profile: "SCHEMATIC1-BIAS"  [ C:\Users\labo\Desktop\402pm\Labo 3 MOS1\ampli source commune-pspicefiles\schematic1\bias.sim ] 

** Creating circuit file "BIAS.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "C:/Users/labo/Desktop/402/Libraries for ELEC-H402/SEDRA_LIB.lib" 
* From [PSPICE NETLIST] section of C:\OrCAD\OrCAD_16.3_Demo\tools\PSpice\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
