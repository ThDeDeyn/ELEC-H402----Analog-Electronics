** Profile: "SCHEMATIC1-Xfert"  [ D:\PM\Documents PM\Cours\_Analogique\ELEC-H-402 2013-2014\Labos\Labo4 MOS2\Ampli Drain Commun\amplidraincommun-pspicefiles\schematic1\xfert.sim ] 

** Creating circuit file "Xfert.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "D:/pm/Documents PM/Cours/_Analogique/ELEC-H-402 2011-2012/Labos/Labo H402 PSpice Lib/small_signal.lib" 
* From [PSPICE NETLIST] section of C:\Program Files\CAO\OrCAD_16.3_Demo\tools\PSpice\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN V_VGQ 0 5 .01 
.STEP PARAM RSval LIST 1u,10 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
